module MY_AND2 (input A,
	     input B,
	     output Z);
assign Z = A & B;
endmodule
